library verilog;
use verilog.vl_types.all;
entity DEUARC_Mesut_Selim_Serbes_2017510100 is
    port(
        outputRegister  : out    vl_logic_vector(3 downto 0);
        Clock           : in     vl_logic;
        InputRegister_in: in     vl_logic_vector(3 downto 0)
    );
end DEUARC_Mesut_Selim_Serbes_2017510100;
