library verilog;
use verilog.vl_types.all;
entity DEUARC_Mesut_Selim_Serbes_2017510100_vlg_vec_tst is
end DEUARC_Mesut_Selim_Serbes_2017510100_vlg_vec_tst;
