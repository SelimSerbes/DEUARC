library verilog;
use verilog.vl_types.all;
entity DEUARC_Mesut_Selim_Serbes_2017510100_vlg_check_tst is
    port(
        outputRegister  : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end DEUARC_Mesut_Selim_Serbes_2017510100_vlg_check_tst;
