library verilog;
use verilog.vl_types.all;
entity DEUARC_Mesut_Selim_Serbes_2017510100_vlg_sample_tst is
    port(
        Clock           : in     vl_logic;
        InputRegister_in: in     vl_logic_vector(3 downto 0);
        sampler_tx      : out    vl_logic
    );
end DEUARC_Mesut_Selim_Serbes_2017510100_vlg_sample_tst;
